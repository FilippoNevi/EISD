library ieee;
use ieee.std_logic_1164.all;

use ieee.upf.all;

entity motor_long_tb is
end entity motor_long_tb;

