`line 4
module vloga_dig_submod_motor_long_tb(\_adms_signal_#dummy\ );
output  \_adms_signal_#dummy\  ;
endmodule

