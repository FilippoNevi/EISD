* Temporary input file

.model motor_long_tb macro lang=veriloga
ytop motor_long_tb

.tran 1u 10sec
//.OPTION HMAX=1u
//.OPTION HMIN=1u
//.ac dec 1k 1 10G
