library ieee;
use ieee.std_logic_1164.all;

use ieee.upf.all;

entity diode_circuit_tb is
end entity diode_circuit_tb;

