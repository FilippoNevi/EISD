LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

LIBRARY STD;
USE STD.ALL;

ENTITY vsrc IS
  PORT (
    SIGNAL p : OUT STD_LOGIC;
    SIGNAL n : OUT STD_LOGIC;
    SIGNAL dc : IN STD_LOGIC_VECTOR(9 downto 0) );
END ENTITY vsrc;

