`line 4
module vloga_dig_submod_diode_circuit_tb(\_adms_signal_#dummy\ );
output  \_adms_signal_#dummy\  ;
endmodule

